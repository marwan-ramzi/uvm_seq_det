`define LENGTH 4
